// Minimal gemm_accelerator.v stub to allow Verilator to build simulation
// This is a simplified stub for simulation purposes only.
module gemm_accelerator (
    input        clk,
    input        rst_n,
    input        start,
    output reg   done,
    output reg   busy,
    // AXI-lite slave signals (simplified)
    input  [31:0] s_axi_awaddr,
    input         s_axi_awvalid,
    output reg    s_axi_awready,
    input  [31:0] s_axi_wdata,
    input  [3:0]  s_axi_wstrb,
    input         s_axi_wvalid,
    output reg    s_axi_wready,
    output reg    s_axi_bvalid,
    input         s_axi_bready
);

    initial begin
        s_axi_awready = 1'b0;
        s_axi_wready  = 1'b0;
        s_axi_bvalid  = 1'b0;
        done = 1'b0;
        busy = 1'b0;
    end

    // Simple behavior: accept writes and return bvalid, respond to start by asserting done next cycle
    always @(posedge clk) begin
        if (!rst_n) begin
            s_axi_awready <= 1'b0;
            s_axi_wready  <= 1'b0;
            s_axi_bvalid  <= 1'b0;
            done <= 1'b0;
            busy <= 1'b0;
        end else begin
            s_axi_awready <= s_axi_awvalid;
            s_axi_wready  <= s_axi_wvalid;
            s_axi_bvalid  <= s_axi_awvalid & s_axi_wvalid;

            if (start) begin
                busy <= 1'b1;
                done <= 1'b0;
            end

            // simulate quick operation: done on next clock
            if (busy) begin
                done <= 1'b1;
                busy <= 1'b0;
            end

            if (s_axi_bvalid && s_axi_bready) begin
                s_axi_bvalid <= 1'b0;
            end
        end
    end
endmodule
// Simple GEMM Accelerator Top Module
// This is a minimal implementation for testing the build system

`timescale 1ns / 1ps

module gemm_accelerator #(
    parameter PE_ROWS = 8,
    parameter PE_COLS = 8,
    parameter DATA_WIDTH = 16,
    parameter ADDR_WIDTH = 32,
    parameter ACC_WIDTH = 32
) (
    input wire clk,
    input wire rst_n,
    
    // AXI4-Lite Configuration Interface (simplified)
    input wire [ADDR_WIDTH-1:0] s_axi_awaddr,
    input wire s_axi_awvalid,
    output reg s_axi_awready,
    input wire [31:0] s_axi_wdata,
    input wire [3:0] s_axi_wstrb,
    input wire s_axi_wvalid,
    output reg s_axi_wready,
    output reg [1:0] s_axi_bresp,
    output reg s_axi_bvalid,
    input wire s_axi_bready,
    
    input wire [ADDR_WIDTH-1:0] s_axi_araddr,
    input wire s_axi_arvalid,
    output reg s_axi_arready,
    output reg [31:0] s_axi_rdata,
    output reg [1:0] s_axi_rresp,
    output reg s_axi_rvalid,
    input wire s_axi_rready,
    
    // Memory Interface - Simplified for testing
    output reg [ADDR_WIDTH-1:0] mem_a_addr,
    output reg mem_a_en,
    input wire [DATA_WIDTH*PE_COLS-1:0] mem_a_data,
    input wire mem_a_valid,
    
    output reg [ADDR_WIDTH-1:0] mem_b_addr,
    output reg mem_b_en,
    input wire [DATA_WIDTH*PE_ROWS-1:0] mem_b_data,
    input wire mem_b_valid,
    
    output reg [ADDR_WIDTH-1:0] mem_c_addr,
    output reg mem_c_en,
    output reg mem_c_we,
    output reg [ACC_WIDTH*PE_ROWS*PE_COLS-1:0] mem_c_data,
    output reg mem_c_valid,
    
    // Status and Control
    output reg busy,
    output reg done,
    input wire start
);

    // Configuration Registers
    reg [15:0] matrix_m, matrix_n, matrix_k;
    reg [1:0] data_format;
    reg accumulate_mode;
    reg [31:0] cycles_counter;
    
    // Control FSM States
    localparam IDLE = 3'b000,
               LOAD = 3'b001,
               COMPUTE = 3'b010,
               STORE = 3'b011,
               DONE = 3'b100;
    
    reg [2:0] state, next_state;
    
    // Initialize registers
    initial begin
        state = IDLE;
        matrix_m = 64;
        matrix_n = 64;
        matrix_k = 64;
        data_format = 2'b10; // INT16
        accumulate_mode = 1'b0;
        cycles_counter = 0;
        busy = 1'b0;
        done = 1'b0;
        
        // Initialize AXI signals
        s_axi_awready = 1'b0;
        s_axi_wready = 1'b0;
        s_axi_bresp = 2'b00;
        s_axi_bvalid = 1'b0;
        s_axi_arready = 1'b0;
        s_axi_rdata = 32'h0;
        s_axi_rresp = 2'b00;
        s_axi_rvalid = 1'b0;
        
        // Initialize memory interface
        mem_a_addr = 0;
        mem_a_en = 1'b0;
        mem_b_addr = 0;
        mem_b_en = 1'b0;
        mem_c_addr = 0;
        mem_c_en = 1'b0;
        mem_c_we = 1'b0;
        mem_c_data = 0;
        mem_c_valid = 1'b0;
    end
    
    // Simple FSM for testing
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            cycles_counter <= 0;
            busy <= 1'b0;
            done <= 1'b0;
        end else begin
            cycles_counter <= cycles_counter + 1;
            
            case (state)
                IDLE: begin
                    busy <= 1'b0;
                    done <= 1'b0;
                    if (start) begin
                        state <= COMPUTE;
                        busy <= 1'b1;
                    end
                end
                
                COMPUTE: begin
                    // Simulate computation time
                    if (cycles_counter > 1000) begin
                        state <= DONE;
                        busy <= 1'b0;
                        done <= 1'b1;
                    end
                end
                
                DONE: begin
                    state <= IDLE;
                    done <= 1'b0;
                    cycles_counter <= 0;
                end
                
                default: state <= IDLE;
            endcase
        end
    end
    
    // Simple AXI4-Lite read interface
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            s_axi_arready <= 1'b0;
            s_axi_rvalid <= 1'b0;
            s_axi_rdata <= 32'h0;
        end else begin
            if (s_axi_arvalid && !s_axi_rvalid) begin
                s_axi_arready <= 1'b1;
                s_axi_rvalid <= 1'b1;
                
                case (s_axi_araddr[7:0])
                    8'h00: s_axi_rdata <= {16'h0, matrix_m};
                    8'h04: s_axi_rdata <= {16'h0, matrix_n};
                    8'h08: s_axi_rdata <= {16'h0, matrix_k};
                    8'h1C: s_axi_rdata <= {30'h0, done, busy};
                    8'h20: s_axi_rdata <= cycles_counter;
                    default: s_axi_rdata <= 32'hDEADBEEF;
                endcase
            end else begin
                s_axi_arready <= 1'b0;
                if (s_axi_rready) begin
                    s_axi_rvalid <= 1'b0;
                end
            end
        end
    end
    
    // Simple AXI4-Lite write interface
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            s_axi_awready <= 1'b0;
            s_axi_wready <= 1'b0;
            s_axi_bvalid <= 1'b0;
        end else begin
            // Simplified write handling
            if (s_axi_awvalid && s_axi_wvalid && !s_axi_bvalid) begin
                s_axi_awready <= 1'b1;
                s_axi_wready <= 1'b1;
                s_axi_bvalid <= 1'b1;
                
                case (s_axi_awaddr[7:0])
                    8'h00: matrix_m <= s_axi_wdata[15:0];
                    8'h04: matrix_n <= s_axi_wdata[15:0];
                    8'h08: matrix_k <= s_axi_wdata[15:0];
                    8'h0C: data_format <= s_axi_wdata[1:0];
                endcase
            end else begin
                s_axi_awready <= 1'b0;
                s_axi_wready <= 1'b0;
                if (s_axi_bready) begin
                    s_axi_bvalid <= 1'b0;
                end
            end
        end
    end

endmodule